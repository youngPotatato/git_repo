class my_env extends uvm_env;
	`uvm_component_utils(my_env)


	function new(string name, uvm_component parent);
		super.new(name,parent);
	endfunction:new

	function void build_phase(uvm_phase phase);
		super.build_phase(phase);
	endfunction:build_phase

	task run_phase(uvm_phase phase);
		phase.raise_object(this);
		#10;
		phase.drop_objection(this);
	endtask:run_phase
endclass:my_env
