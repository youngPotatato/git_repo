
// DEFINES 
`define __FILE__ "NA.v"
`define __LINE__ 0
`define __VAMS_ENABLE__
`define __VAMS_COMPACT_MODELING__
`define DVT_PATCH

// CONFIGURATION FILES (libmap) 
`include "/home/yy/EDA/uvm-1.2/src/uvm_pkg.sv"
`include "/home/yy/Desktop/My_prog/git_repo/DVT_PROJ/1/uvm-1.2_ubus/examples/ubus_tb_top.sv"
