`timescale 1ns/1ns
parameter cycle = 100;	
typedef enum {ADD,SUB,MULT,DIV} opcode_e;

