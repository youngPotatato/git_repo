`define Width 16 
`define Depth_bits 7 
