typedef uvm_sequencer #(my_transaction_base) my_sequencer;
