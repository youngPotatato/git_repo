
// DEFINES 
`define __FILE__ "NA.v"
`define __LINE__ 0
`define __VAMS_ENABLE__
`define __VAMS_COMPACT_MODELING__
`define DVT_PATCH

// CONFIGURATION FILES (libmap) 
`include "/home/yy/Desktop/My_prog/git_repo/DVT_PROJ/1/sv-GettingStarted/defines.sv"
`include "/home/yy/Desktop/My_prog/git_repo/DVT_PROJ/1/sv-GettingStarted/class_1.sv"
`include "/home/yy/Desktop/My_prog/git_repo/DVT_PROJ/1/sv-GettingStarted/class_2.sv"
`include "/home/yy/Desktop/My_prog/git_repo/DVT_PROJ/1/sv-GettingStarted/class_3.sv"
`include "/home/yy/Desktop/My_prog/git_repo/DVT_PROJ/1/sv-GettingStarted/class_4.sv"
`include "/home/yy/Desktop/My_prog/git_repo/DVT_PROJ/1/sv-GettingStarted/class_5.sv"
