`define Width 16 
`define Depth_bits 2 
`define Max_Ratio 16// the ratio of Max randomized trasa num over 
		    // the depth of lifo/fifo
