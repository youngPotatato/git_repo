`ifndef ENV_SVH
`define ENV_SVH

import uvm_pkg::*;

`include "uvm_macros.svh"
`include "../test/definition.sv"
`include "../test/dut_if.sv"
`include "transfer.sv"
`include "my_sequencer.sv"
`include "my_dut_config.sv"
`include "my_driver.sv"
`include "my_monitor.sv"
`include "my_agent.sv"
`include "my_scoreboard.sv"
`include "my_env.sv"


`endif // ENV_SVH
