module dut(dut_if _if); 
	always @(posedge _if.clk) begin
	end
endmodule:dut
