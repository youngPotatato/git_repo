

class class_4 extends class_2;

    // HINT Learn about rename refactoring
    //
    // Click 'too' and
    //   right-click to Refactor > Rename
    //   or press Alt+Shift+R
    //
    // to rename 'too' into 'tootoo'.
    //
    // Preview changes across all relevant files and press OK in the dialog to rename.
    //
    // Note that 'v5.too()' below is not changed.
    //
    // Rename works for any identifier (variables, functions, classes, macros etc.).
    virtual task too();
        class_5 v5;

        super.too();

        v5.too();
    endtask


    // HINT Learn about Override Methods Wizard
    //
    // Type 'foo', press Ctrl+Space, chose Override Methods..., and press Enter.
    //
    // Once you override the method you should get something like:
    //
    // virtual function int foo_1();
    //     // TODO Auto-generated function stub
    //     return super.foo_1();
    // endfunction : foo_1


    // HINT Learn about code formatting
    //
    // If the source code is not properly aligned:
    //   right-click in the editor and Source > Format Source
    //   or press Ctrl+Shift+F


    // HINT Learn about hyperlinks
    //
    // Ctrl+click 'fld5' to open field type.
    local class_5 fld5;

endclass
