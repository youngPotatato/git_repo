interface dut_if();
endinterface:dut_if
