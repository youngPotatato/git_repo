interface dut_if;
	lobic rst,clk;
	logic data;
endinterface:dut_if
