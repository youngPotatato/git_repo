
// DEFINES 
`define __FILE__ "NA.v"
`define __LINE__ 0
`define __VAMS_ENABLE__
`define __VAMS_COMPACT_MODELING__
`define DVT_PATCH
`define LITLE_ENDIAN
`define UART_ABV_ON
`define INCA
`define wrealXState 0
`define wrealZState 0

// CONFIGURATION FILES (libmap) 
`include "/home/yy/EDA/dvt_eclipse/predefined_projects/libs/uvm-1.1b/src/uvm_pkg.sv"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/opencores/uart16550/rtl/uart_defines.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/opencores/spi/rtl/spi_defines.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/soc_verification_lib/sv_cb_ex_lib/apb_subsystem/sv/gpio_defines.svh"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/soc_verification_lib/sv_cb_ex_lib/apb_subsystem/sv/spi_defines.svh"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/soc_verification_lib/sv_cb_ex_lib/uart_ctrl/sv/uart_ctrl_defines.svh"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/soc_verification_lib/sv_cb_ex_lib/apb_subsystem/sv/apb_subsystem_defines.svh"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/soc_verification_lib/sv_cb_ex_lib/interface_uvc_lib/ahb/sv/ahb_pkg.sv"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/soc_verification_lib/sv_cb_ex_lib/interface_uvc_lib/apb/sv/apb_pkg.sv"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/soc_verification_lib/sv_cb_ex_lib/interface_uvc_lib/uart/sv/uart_pkg.sv"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/soc_verification_lib/sv_cb_ex_lib/interface_uvc_lib/gpio/sv/gpio_pkg.sv"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/soc_verification_lib/sv_cb_ex_lib/interface_uvc_lib/spi/sv/spi_pkg.sv"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/soc_verification_lib/sv_cb_ex_lib/uart_ctrl/sv/uart_ctrl_pkg.sv"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/soc_verification_lib/sv_cb_ex_lib/apb_subsystem/sv/apb_subsystem_pkg.sv"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/soc_verification_lib/sv_cb_ex_lib/apb_subsystem/tb/sv/apb_subsystem_top.sv"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/apb_subsystem/rtl/apb_subsystem_0.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/apb_subsystem/rtl/apb_subsystem_1.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/apb_subsystem/rtl/alut_veneer.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/apb_subsystem/rtl/gpio_veneer.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/apb_subsystem/rtl/ttc_veneer.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/apb_subsystem/rtl/smc_veneer.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/apb_subsystem/rtl/power_ctrl_veneer.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/ahb2apb/rtl/ahb2apb.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/alut/rtl/alut_reg_bank.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/alut/rtl/alut_addr_checker.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/alut/rtl/alut_mem.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/alut/rtl/alut_age_checker.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/alut/rtl/alut.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/opencores/spi/rtl/spi_clgen.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/opencores/spi/rtl/spi_shift.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/opencores/spi/rtl/spi_top.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/opencores/uart16550/rtl/uart_top.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/opencores/uart16550/rtl/uart_wb.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/opencores/uart16550/rtl/uart_transmitter.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/opencores/uart16550/rtl/uart_receiver.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/opencores/uart16550/rtl/uart_tfifo.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/opencores/uart16550/rtl/uart_rfifo.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/opencores/uart16550/rtl/uart_regs.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/opencores/uart16550/rtl/uart_debug_if.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/opencores/uart16550/rtl/raminfr.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/opencores/uart16550/rtl/uart_sync_flops.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/gpio/rtl/gpio_lite_subunit.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/gpio/rtl/gpio_lite.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/ttc/rtl/ttc_counter_lite.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/ttc/rtl/ttc_interface_lite.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/ttc/rtl/ttc_interrupt_lite.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/ttc/rtl/ttc_count_rst_lite.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/ttc/rtl/ttc_timer_counter_lite.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/ttc/rtl/ttc_lite.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/smc/rtl/smc_addr_lite.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/smc/rtl/smc_cfreg_lite.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/smc/rtl/smc_apb_lite_if.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/smc/rtl/smc_ahb_lite_if.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/smc/rtl/smc_counter_lite.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/smc/rtl/smc_mac_lite.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/smc/rtl/smc_state_lite.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/smc/rtl/smc_strobe_lite.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/smc/rtl/smc_wr_enable_lite.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/smc/rtl/smc_lite.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/power_ctrl/rtl/power_ctrl_sm.v"
`include "/home/yy/dvt_predefined_projects_target/uvm_ref_flow_1.1/designs/socv/rtl/rtl_lpw/power_ctrl/rtl/power_ctrl.v"
