module dut(dut_if _if);
endmodule:dut
