package my_pkg;
	`include "uvm_macros.svh"
	import uvm_pkg::*;
	`include "environment.sv"
	`include "test.sv"
endpackage:my_pkg
